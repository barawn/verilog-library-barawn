`timescale 1ns / 1ps
`include "dsp_macros.vh"

// (C) Patrick Allison (allison.122@osu.edu) or the Ohio State University.
// Please contact me either directly or via GitHub for reuse purposes.

// This is the compensating FIR for a biquad's pole pair.
// v2 rearranges things to reduce power consumption by sharing delays
// and passing the delayed inputs along for the incremental version.
//
// There are two compensating FIRs, one for each of the samples
// generated from the IIR. Sample 0's FIR is called the f chain,
// and sample 1's FIR is called the g chain. These compensating FIRs
// are then pipelined to generate the F and G outputs. One of those
// DSPs is at the end of each of the f/g chains, and then the second
// set of DSPs, which links the two chains, are separate.
//
// The total F chain (consisting of the f and the final pipeline DSP)
// is NSAMP-1 DSPs long.
// The total G chain (consisting of the g and the final pipeline DSP)
// is NSAMP DSPs long.
//
// Because of the difference in total length, the delays between the
// inputs of the two chains differ. The f chain wants to take in
// x[0], x[NSAMP-1]z^-1, x[NSAMP-2]z^-1 ... x[2]z^-1
// and the g chain wants to take in
// x[1], x[0], x[NSAMP-1]z^-1, x[NSAMP-2]z^-1 ... x[2]z^-1
//
// The first dspA output gives (c*x[0]z^-1 + x[1]z^-1)z^-1 or
// c*x[0]z^-2 + x[1]z^-2.
// etc.
// For the most part this is straightforward, we just need to handle the G chain head
// differently.
//
// F chain:     (-P^M)*U_(M-2)(cos t)
//              P*U_1(cos t) ..             (coeff for x[M-2])
//              P^(M-2)U_(M-2)(cos t)       (coeff for x[2])
// G chain:     P^M*U_M(cos t)
//              P^2 U_(M-2)(cos t)          (coeff for x[M-1])
//              ...
//              P^(M-1)U_(M-1)(cos t)       (coeff for x[2])
//              P*U_1(cos t)                (coeff for x[0])
module biquad8_pole_fir_v2 #(parameter NBITS=16, 
                          parameter NFRAC=2,
                          parameter CLKTYPE="NONE",
                          parameter NSAMP=8,
                          // How many clocks after 'bypass_i' changes
                          // do we expect bypassed/unbypassed data
                          // to show up.
                          parameter BYPASS_DELAY=3) (
        input			clk,
        input [NBITS*NSAMP-1:0]	dat_i,

        // The bypass input forces all of the MREGs to zero sequentially,
        // converting "y0_out" = sample 0 and "y1_out" = sample 1.
        
        input           bypass_i,
        output          bypass_o,

        // the address here selects
        // 00 : F chain
        // 01 : G chain
        // 10 : F cross-link
        // 11 : G cross-link
        input [1:0]		coeff_adr_i, 
        input			coeff_wr_i,
        input			coeff_update_i,
        input [17:0]		coeff_dat_i,
                
        output [47:0]		y0_out,
        output [47:0]		y1_out,
        // Delayed versions of the input, with increasing delays.
        // Each input past 2 has (sample-2) clocks of delay.
        output [NBITS*NSAMP-1:0] x_out
    );

    // Total length of the F chain = (f length + 1)
    localparam FLEN = NSAMP-1;
    // Total length of the G chain = (g length + 1)
    localparam GLEN = NSAMP;
    
    // Outputs and cascades from the F chain    
    wire [47:0] fpout[FLEN-1:0];
    wire [17:0] fbcascade[FLEN-1:0];
    wire [47:0] fpcascade[FLEN-1:0];
    // Outputs and cascades from the G chain
    wire [17:0] gbcascade[GLEN-1:0];
    wire [47:0] gpcascade[GLEN-1:0];
    wire [47:0] gpout[GLEN-1:0];
    
    // after bypass, there are BYPASS_DELAY clocks before bypassed
    // data starts showing up.
    wire [FLEN-1:0] force_f_bypass;
    wire [GLEN-1:0] force_g_bypass;
    // g chain delays RSTM by BYPASS_DELAY+1 clocks, f chain delays
    // by BYPASS_DELAY+2 clocks.
    reg [BYPASS_DELAY+1:0] bypass_shreg = {(BYPASS_DELAY+2){1'b0}};

    wire f_bypass_in = bypass_shreg[BYPASS_DELAY+1];
    wire g_bypass_in = bypass_shreg[BYPASS_DELAY];

    // Registered control signals.
    (* CUSTOM_CC_DST = CLKTYPE *)
    reg coeff_wr_f = 0;
    (* CUSTOM_CC_DST = CLKTYPE *)
    reg coeff_wr_g = 0;
    (* CUSTOM_CC_DST = CLKTYPE *)
    reg	coeff_wr_fcross = 0;
    (* CUSTOM_CC_DST = CLKTYPE *)
    reg	coeff_wr_gcross = 0;   
  
    // Update all coefficients.
    reg update = 0;

    // Logic for coefficient control.
    integer b;
    always @(posedge clk) begin
       for (b=0;b<(BYPASS_DELAY+2);b=b+1) begin
           bypass_shreg[b] <= (b==0) ? bypass_i : bypass_shreg[b-1];
       end
       coeff_wr_f <= coeff_wr_i && (coeff_adr_i == 2'b00);       
       coeff_wr_g <= coeff_wr_i && (coeff_adr_i == 2'b01);

       update <= coeff_update_i;

       coeff_wr_fcross <= coeff_wr_i && (coeff_adr_i == 2'b10);
       coeff_wr_gcross <= coeff_wr_i && (coeff_adr_i == 2'b11);       
    end

    `define COMMON_ATTRS    `CONSTANT_MODE_ATTRS, `DE2_UNUSED_ATTRS, .BREG(2), .BCASCREG(1), .PREG(1)    

    // Our goal here is to allow as many registers here to be shared as
    // possible. Looking at NSAMP=4 and assuming AREG=1, MREG=1, CREG=1, that means
    // the PREG output is delayed 3 clocks.
    // A -> z^-1 (AREG)    z^-1(MREG)       \
    // C -> z^-1 (CREG)                     +-- z^-1 (PREG) ==>
    //
    // e.g. P output = (B*Az^-2 + Cz^-1)z^-1
    //
    // Considering the g chain first because it's longer:
    // dspA's P output: (BA*x[0]z^-2 + C(x[1]z^-1)z^-1)z^-1 = dspA at z^-3
    // dspB's P output: (BB*(x[2]z^-1)z^-2 + dspA)z^-1 = dspB at z^-4
    // dspC's P output: (BC*(x[3]z^-2)z^-2 + dspB)z^-1 = dspC at z^-5
    //
    // Now the f chain needs:
    // dspA's P output: (BA*(x[2]z^-1)z^-2 + C(x[0]z^-2)z^-1)z^-1 = dspA at z^-4
    // dspB's P output: (BB*(x[3]z^-2)z^-2 + dspA)z^-1 = dspB at z^-5
    //
    // This means we need:
    // x[0] and x[0]z^-2
    // x[1]z^-1
    // x[2]z^-1
    // x[3]z^-2
    // etc.
    //
    // BYPASS_DELAY is the amount of time from bypass_i until
    // bypassed data shows up at the input. e.g. if BYPASS_DELAY=3,
    // and bypass turns on at clock 1, it shows up at clock 4.
    // For the f-chain, we want
    //
    // clk  bypass  RSTM    FIR2    A           AREG        MREG            C           CREG        PREG
    // 0    0       0       FIR2[0] FIR2[-1]    FIR2[-2]    BA*FIR2[-3]     FIR0[-2]    FIR0[-3]    FIR0[-4]+BA*FIR2[-4]
    // 1    1       0       FIR2[1] FIR2[0]     FIR2[-1]    BA*FIR2[-2]     FIR0[-1]    FIR0[-2]    FIR0[-3]+BA*FIR2[-3]
    // 2    1       0       FIR2[2] FIR2[1]     FIR2[0]     BA*FIR2[-1]     FIR0[0]     FIR0[-1]    FIR0[-2]+BA*FIR2[-2]
    // 3    1       0       FIR2[3] FIR2[2]     FIR2[1]     BA*FIR2[0]      FIR0[1]     FIR0[0]     FIR0[-1]+BA*FIR2[-1]
    // 4    1       0       D[4]    FIR2[3]     FIR2[2]     BA*FIR2[1]      FIR0[2]     FIR0[1]     FIR0[0]+BA*FIR2[0]
    // 5    1       0       D[5]    D[4]        FIR2[3]     BA*FIR2[2]      FIR0[3]     FIR0[2]     FIR0[1]+BA*FIR2[1]
    // 6    1       1       D[6]    D[5]        D[4]        BA*FIR2[3]      D[4]        FIR0[3]     FIR0[2]+BA*FIR2[2]
    // 7    1       1       D[7]    D[6]        D[5]        0               D[5]        D[4]        FIR0[3]+BA*FIR2[3]
    // 8    1       1       D[8]    D[7]        D[6]        0               D[6]        D[5]        D[4]
    // which means the F-chain's first RSTM is the output of a 5 clock shift reg
    // dspA RSTM = bypass_shreg[4]
    // dspB RSTM = bypass_shreg[5]
    // dspC RSTM = bypass_shreg[6]
    //
    // The g-chain is one shorter:
    // 
    // clk  bypass  RSTM    FIR0    A           AREG        MREG            C           CREG        PREG
    // 0    0       0       FIR0[0] FIR0[0]     FIR0[-1]    BA*FIR0[-2]     FIR1[-1]    FIR1[-2]    FIR1[-3]+BA*FIR0[-3]
    // 1    1       0       FIR0[1] FIR0[1]     FIR0[0]     BA*FIR0[-1]     FIR0[0]     FIR1[-1]    FIR1[-2]+BA*FIR0[-2]
    // 2    1       0       FIR0[2] FIR0[2]     FIR0[1]     BA*FIR0[0]      FIR0[1]     FIR1[0]     FIR1[-1]+BA*FIR0[-1]
    // 3    1       0       FIR0[3] FIR0[3]     FIR0[2]     BA*FIR0[1]      FIR0[2]     FIR1[1]     FIR1[0]+BA*FIR0[0]
    // 4    1       0       D[4]    D[4]        FIR0[3]     BA*FIR0[2]      FIR0[3]     FIR1[2]     FIR1[1]+BA*FIR0[1]
    // 5    1       1       D[5]    D[5]        D[4]        BA*FIR0[3]      D[4]        FIR1[3]     FIR1[2]+BA*FIR0[2]
    // 6    1       1       D[6]    D[6]        D[5]        0               D[5]        D[4]        FIR1[3]+BA*FIR0[3]
    // 7    1       1       D[7]    D[7]        D[6]        0               D[6]        D[5]        D[4]
    
    // so for the g chain
    // dspA RSTM = bypass_shreg[3]  turns on at clk7 after clk1
    // dspB RSTM = bypass_shreg[4]  turns on at clk8 after clk1
    // dspC RSTM = bypass_shreg[5]  turns on at clk9 after clk1
    // dspD RSTM = bypass_shreg[6]  turns on at clk10 after clk1
    // 
        
    // The g chain is NSAMP clocks long:
    //
    // 
    //
    // f        dspA ALU in             dspA P      dspB
    // x[0]     x[0][-3] + B*x[2][-3]
    // x[2]     
    // x[3]                             x[0][-4] + B*x[2][-4] + C*x[3][-4]

    // So clearly x[1] needs a delay of 1 clock

    // g        dspA                    dspB                        dspC
    // x[1]     x[1][-2] + D*x[0][-2]
    // x[0]
    // x[2]                             x[1][-3]+Dx[0][-3]+Ex[2][-3]
    // x[3]                                                         x[1][-4]+Dx[0][-4]+Ex[2][-4]+Fx[3][-4]
    // CHEAP IMPROVEMENT
    // What we were PREVIOUSLY doing was 
    // 7    -> SRL(A=2)->FF ->  F dspA_in[0]
    //      -> SRL(A=1)->FF ->  G dspA_in[1]
    // 6    -> SRL(A=3)->FF ->  F dspA_in[1]
    //      -> SRL(A=2)->FF ->  G dspA_in[2]
    // etc.
    // This is obviously dumb. We can just do
    // 7    -> SRL(A=1)->FF ->  G dspA_in[1]
    //                   |--->  F dspA_in[0] with an extra AREG.
    //
    // Additionally, there's no reason for us to arrange the chains in any particular order at all.
    // Note that here, we end up with sample 7 with the shortest delays,
    // then sample 6, then sample 5, etc.
    // But for the incremental computation portion, sample 7 will end up needing the longest delay.
    // So instead, reverse this. It's just a change of programming parameters. And then actually
    // output all of the delayed values so we can reuse them in the incremental without
    // adding more delays.
    
    wire [NSAMP-1:0][NBITS-1:0] in_delayed;  
    
    localparam NUM_HEAD_PAD = 17 - (NBITS-NFRAC);
    localparam NUM_TAIL_PAD = 13 - NFRAC;

    generate    
        genvar fi,fj, gi,gj, smp;

        // Generate the delays.
        for (smp=0;smp<NSAMP;smp=smp+1) begin : DLY
            // sample 0 gets 2 clocks, sample 1 gets 1 clock,
            // sample 2 gets 2 clocks
            // sample 3 gets 3 clocks
            // sample 4 gets 4 clocks, etc.
            localparam DELAY = (smp < 2) ? ((smp < 1) ? 2 : 1) : (2 + (smp-2));
            reg [DELAY-1:0][NBITS-1:0] in_store = {NBITS*DELAY{1'b0}};
            integer s;
            always @(posedge clk) begin : ST
                for (s=0;s<DELAY;s=s+1) begin : LP
                    in_store[s] <= (s==0) ? dat_i[NBITS*smp +: NBITS] : in_store[s-1];
                end
            end
            assign in_delayed[smp] = in_store[DELAY-1];
            assign x_out[NBITS*smp +: NBITS] = in_delayed[smp];
        end
        // Now run the f chain.        
        for (fi=0;fi<FLEN;fi=fi+1) begin : FLOOP
            reg rstm = 0;
            always @(posedge clk) begin : RB
                rstm <= (fi == 0) ? f_bypass_in : force_f_bypass[fi-1];
            end
            assign force_f_bypass[fi] = rstm;
            // F chain has AREG=2-FABRIC_DELAY, ADREG=0, MREG=1
            wire [29:0] dspA_in = (fi < FLEN-1) ?
                { {NUM_HEAD_PAD{in_delayed[fi+2][NBITS-1]}}, in_delayed[fi+2], {NUM_TAIL_PAD{1'b0}} } :
                  fpout[fi-1][14 +: 30];

            if (fi == 0) begin : HEAD
                localparam THIS_AREG = 1;
                wire THIS_CEA1 = (THIS_AREG > 1) ? 1'b1 : 1'b0;
                wire THIS_CEA2 = (THIS_AREG > 0) ? 1'b1 : 1'b0;
                localparam C_HEAD_PAD = 21 - (NBITS-NFRAC);
                localparam C_TAIL_PAD = 27 - NFRAC;
                // in_delayed[0] is delayed by 2 clocks.
                wire [47:0] dspC_in = { {C_HEAD_PAD{in_delayed[0][NBITS-1]}}, in_delayed[0], {C_TAIL_PAD{1'b0}} };
                // the f chain will have AREG=2, ADREG=0, MREG=1                
                (* CUSTOM_CC_DST = CLKTYPE *)
                DSP48E2 #(`COMMON_ATTRS,
                          .CREG(1),
                          .AREG(THIS_AREG),
                          .ACASCREG(THIS_AREG),
                          .ADREG(0),
                          .MREG(1))
                    u_head( .CLK(clk),
                            .CEP(1'b1),
                            .CEC(1'b1),
                            .CEM(1'b1),
                            .RSTM(rstm),
                            .CEA1(THIS_CEA1),
                            .CEA2(THIS_CEA2),
                            .C(dspC_in),   // This is where the 1 in [1,X_1,X_2,...] is added             
                            .A(dspA_in),
                            .B(coeff_dat_i),
                            .BCOUT(fbcascade[fi]),
                            .CEB1(coeff_wr_f),  // The first clock enable allows the new coefficients to flow in (but not apply)
                            .CEB2(update),      // The second clock eneable applies the coefficients
                            `D_UNUSED_PORTS,
                            .CARRYINSEL(`CARRYINSEL_CARRYIN),
                            .ALUMODE(`ALUMODE_SUM_ZXYCIN),
                            .OPMODE( { 2'b00, `Z_OPMODE_C, `XY_OPMODE_M } ),
                            .INMODE( 0 ),
                            .P(fpout[fi]),
                            .PCOUT(fpcascade[fi]));
            end else begin : BODY
                localparam THIS_AREG = (fi < FLEN-1) ? 1 : 0;
                wire THIS_CEA1 = 0;
                wire THIS_CEA2 = (fi < FLEN-1 && THIS_AREG > 0) ? 1 : 0;
                DSP48E2 #(`COMMON_ATTRS,
                          `C_UNUSED_ATTRS,
                          .B_INPUT("CASCADE"),
                          .AREG(THIS_AREG),
                          .ACASCREG(THIS_AREG),
                          .ADREG(0),
                          .MREG(1))
                    u_body( .CLK(clk),
                            .CEP(1'b1),                            
                            .A(dspA_in),
                            .CEA2(THIS_CEA2),
                            .CEA1(THIS_CEA1),
                            .CEM(1'b1),
                            .RSTM(rstm),
                            .BCIN(fbcascade[fi-1]),
                            .BCOUT(fbcascade[fi]),
                            .CEB1(coeff_wr_f),
                            .CEB2(update),
                            `C_UNUSED_PORTS,
                            `D_UNUSED_PORTS,
                            .CARRYINSEL(`CARRYINSEL_CARRYIN),
                            .ALUMODE(`ALUMODE_SUM_ZXYCIN),
                            .OPMODE( { 2'b00, `Z_OPMODE_PCIN, `XY_OPMODE_M } ),
                            .INMODE( 0 ),
                            .P(fpout[fi]),
                            .PCIN(fpcascade[fi-1]),
                            .PCOUT(fpcascade[fi]) );
            end 
        end
        // And the g chain
        for (gi=0;gi<GLEN;gi=gi+1) begin : GLOOP
            reg rstm = 0;
            always @(posedge clk) begin : RB
                rstm <= (gi == 0) ? g_bypass_in : force_g_bypass[gi-1];
            end
            assign force_g_bypass[gi] = rstm;
            localparam int IDX = (gi > 0) ? gi+1 : 0;            
            // g chain's head input is different.

            // head gets AREG=1, MREG=0
            if (gi == 0) begin : HEAD
                localparam C_HEAD_PAD = 21 - (NBITS-NFRAC);
                localparam C_TAIL_PAD = 27 - NFRAC;
                // Head DSP gets x[0] and x[1]z^-1.
                wire [NBITS-1:0] head_input = dat_i[0 +: NBITS];
                wire [29:0] dspA_in = { {NUM_HEAD_PAD{head_input[NBITS-1]}}, head_input, {NUM_TAIL_PAD{1'b0}} };
                wire [47:0] dspC_in = { {C_HEAD_PAD{in_delayed[1][NBITS-1]}}, in_delayed[1], {C_TAIL_PAD{1'b0}} }; 
                // HEAD dsp gets its inputs directly
                (* CUSTOM_CC_DST = CLKTYPE *)
                DSP48E2 #(`COMMON_ATTRS,
                          .CREG(1),
                          .AREG(1),
                          .ADREG(0),
                          .ACASCREG(1),
                          .MREG(1))                          
                    u_head( .CLK(clk),
                            .CEP(1'b1),
                            .CEA2(1'b1),
                            .CEC(1'b1),
                            .CEM(1'b1),
                            .RSTM(rstm),
                            .C(dspC_in),                            
                            .A(dspA_in),
                            .B(coeff_dat_i),
                            .BCOUT(gbcascade[gi]),
                            .CEB1(coeff_wr_g),
                            .CEB2(update),
                            `D_UNUSED_PORTS,
                            .CARRYINSEL(`CARRYINSEL_CARRYIN),
                            .ALUMODE(`ALUMODE_SUM_ZXYCIN),
                            .OPMODE( { 2'b00, `Z_OPMODE_C, `XY_OPMODE_M } ),
                            .INMODE( 0 ),
                            .P(gpout[gi]),
                            .PCOUT(gpcascade[gi]));
            end else begin : BODY
                wire [29:0] dspA_in;
                assign dspA_in = (gi < GLEN-1) ? 
                    { {NUM_HEAD_PAD{in_delayed[IDX][NBITS-1]}}, in_delayed[IDX], {NUM_TAIL_PAD{1'b0}} } :
                      gpout[gi-1][14 +: 30];    
                // and everywhere else gets AREG=2, MREG=1 except the loopback which gets AREG=0           
                localparam THIS_AREG = (gi < GLEN-1) ? 1 : 0;
                wire THIS_CEA1 = 0;
                wire THIS_CEA2 = (gi < GLEN-1 && THIS_AREG > 0) ? 1 : 0;
                DSP48E2 #(`COMMON_ATTRS,
                          .AREG(THIS_AREG),
                          .ACASCREG(THIS_AREG),
                          .MREG(1),
                          .B_INPUT("CASCADE"),
                          `C_UNUSED_ATTRS)
                    u_body( .CLK(clk),
                            .CEP(1'b1),
                            .CEA1(THIS_CEA1),
                            .CEA2(THIS_CEA2),
                            .CEM(1'b1),
                            .RSTM(rstm),
                            .A(dspA_in),
                            .BCIN(gbcascade[gi-1]),
                            .BCOUT(gbcascade[gi]),
                            .CEB1(coeff_wr_g),
                            .CEB2(update),
                            `C_UNUSED_PORTS,
                            `D_UNUSED_PORTS,
                            .CARRYINSEL(`CARRYINSEL_CARRYIN),
                            .ALUMODE(`ALUMODE_SUM_ZXYCIN),
                            .OPMODE( { 2'b00, `Z_OPMODE_PCIN, `XY_OPMODE_M } ),
                            .INMODE( 0 ),
                            .P(gpout[gi]),
                            .PCIN(gpcascade[gi-1]),
                            .PCOUT(gpcascade[gi]) );
            end 
        end
    endgenerate                            
    // Now our final two cross-linked DSPs take fpout[FLEN-2] (=f[n]) and fpout[FLEN-1] = (f[n-1] + B*f[n-2]).
    //
    // We ** might ** want to actually put dspF at the end of the G chain and dspG at the end of the F chain.
    // Right now for instance both GLOOP[7] and dspF both take the same inputs with delay, so there's no reason
    // we couldn't cascade the input there.
    //     
    // plus the equivalent from the G-chain.
    // We want B2*g[n-1] + f[n] + B*f[n-1].
    // So we drop fpout[FLEN-1] into C (meaning it contains f[n-2] and B*f[n-3])
    // and drop gpout[GLEN-2] into A with 2 regs + MREG, meaning
    // A1 contains g[n-1]
    // A2 contains g[n-2]
    // MREG contains B*g[n-3]
    // and equivalent.

    // Grab the bypass from the g chain. Doesn't matter which one.
    // The extra AREG doesn't matter - what matters is at the ALU,
    // since we are computing CREG + MREG. We want to force MREG=0
    // when CREG becomes bypassed, which is one clock after.
    wire cross_bypass_in = force_g_bypass[GLEN-1];
    
    reg cross_bypass = 0;
    reg bypass_output = 0;      
    wire ceb1_f = coeff_wr_fcross;
    wire ceb1_g = coeff_wr_gcross;
    (* KEEP = "TRUE" *)
    reg ceb2_f = 0;
    (* KEEP = "TRUE" *)
    reg ceb2_g = 0;
    always @(posedge clk) begin
        cross_bypass <= cross_bypass_in;
        bypass_output <= cross_bypass;
        ceb2_f <= coeff_update_i;
        ceb2_g <= coeff_update_i;
    end
    // A gets gpout[GLEN-2]
    localparam C_FRAC_BITS = 27;
    localparam A_FRAC_BITS = 13;
    // Then to find where A starts, you just subtract the difference between
    // the A and C frac bits (if they were the same, you start at the same one).
    // Here we drop the bottom 14 bits.
    wire [29:0] dspF_A = { gpout[GLEN-2][(C_FRAC_BITS-A_FRAC_BITS) +: 30] };
    wire [47:0] dspF_C = fpout[FLEN-1];
    (* CUSTOM_CC_DST = CLKTYPE *)
    DSP48E2 #(.AREG(2),.MREG(1),.BREG(2),.PREG(1),.CREG(1),`CONSTANT_MODE_ATTRS,`DE2_UNUSED_ATTRS)
        u_fdsp( .CLK(clk),
                .CEP(1'b1),
                .CEC(1'b1),
                .CEA1(1'b1),
                .CEA2(1'b1),
                .CEM(1'b1),
                .RSTM(cross_bypass),
                .CEB1(ceb1_f),
                .CEB2(ceb2_f),
                .B(coeff_dat_i),
                .A(dspF_A),
                .C(dspF_C),
                .CARRYINSEL(`CARRYINSEL_CARRYIN),
                .ALUMODE(`ALUMODE_SUM_ZXYCIN),
                .OPMODE( { 2'b00, `Z_OPMODE_C, `XY_OPMODE_M } ),
                .INMODE(0),
                .P(y0_out));
    // A gets fpout[GLEN-2]
    wire [29:0] dspG_A = { fpout[FLEN-2][(C_FRAC_BITS-A_FRAC_BITS) +: 30] };
    wire [47:0] dspG_C = gpout[GLEN-1];
    (* CUSTOM_CC_DST = CLKTYPE *)
    DSP48E2 #(.AREG(2),.MREG(1),.BREG(2),.PREG(1),.CREG(1),`CONSTANT_MODE_ATTRS,`DE2_UNUSED_ATTRS)
        u_gdsp( .CLK(clk),
                .CEP(1'b1),
                .CEC(1'b1),
                .CEA1(1'b1),
                .CEA2(1'b1),
                .CEM(1'b1),
                .RSTM(cross_bypass),
                .CEB1(ceb1_g),
                .CEB2(ceb2_g),
                .B(coeff_dat_i),
                .A(dspG_A),
                .C(dspG_C),
                .CARRYINSEL(`CARRYINSEL_CARRYIN),
                .ALUMODE(`ALUMODE_SUM_ZXYCIN),
                .OPMODE( { 2'b00, `Z_OPMODE_C, `XY_OPMODE_M } ),
                .INMODE(0),
                .P(y1_out));

    assign bypass_o = bypass_output;
    
    `undef COMMON_ATTRS
endmodule

